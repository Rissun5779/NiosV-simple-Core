
module Nios_V (
	clk_clk);	

	input		clk_clk;
endmodule
