// Nios_V.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module Nios_V (
		input  wire  clk_clk  // clk.clk
	);

	wire         nios_v_dbg_reset_out_reset;                            // Nios_V:dbg_reset_out_reset -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire  [31:0] nios_v_data_manager_awaddr;                            // Nios_V:data_manager_awaddr -> mm_interconnect_0:Nios_V_data_manager_awaddr
	wire   [1:0] nios_v_data_manager_bresp;                             // mm_interconnect_0:Nios_V_data_manager_bresp -> Nios_V:data_manager_bresp
	wire         nios_v_data_manager_arready;                           // mm_interconnect_0:Nios_V_data_manager_arready -> Nios_V:data_manager_arready
	wire  [31:0] nios_v_data_manager_rdata;                             // mm_interconnect_0:Nios_V_data_manager_rdata -> Nios_V:data_manager_rdata
	wire   [3:0] nios_v_data_manager_wstrb;                             // Nios_V:data_manager_wstrb -> mm_interconnect_0:Nios_V_data_manager_wstrb
	wire         nios_v_data_manager_wready;                            // mm_interconnect_0:Nios_V_data_manager_wready -> Nios_V:data_manager_wready
	wire         nios_v_data_manager_awready;                           // mm_interconnect_0:Nios_V_data_manager_awready -> Nios_V:data_manager_awready
	wire         nios_v_data_manager_rready;                            // Nios_V:data_manager_rready -> mm_interconnect_0:Nios_V_data_manager_rready
	wire         nios_v_data_manager_bready;                            // Nios_V:data_manager_bready -> mm_interconnect_0:Nios_V_data_manager_bready
	wire         nios_v_data_manager_wvalid;                            // Nios_V:data_manager_wvalid -> mm_interconnect_0:Nios_V_data_manager_wvalid
	wire  [31:0] nios_v_data_manager_araddr;                            // Nios_V:data_manager_araddr -> mm_interconnect_0:Nios_V_data_manager_araddr
	wire   [2:0] nios_v_data_manager_arprot;                            // Nios_V:data_manager_arprot -> mm_interconnect_0:Nios_V_data_manager_arprot
	wire   [1:0] nios_v_data_manager_rresp;                             // mm_interconnect_0:Nios_V_data_manager_rresp -> Nios_V:data_manager_rresp
	wire   [2:0] nios_v_data_manager_awprot;                            // Nios_V:data_manager_awprot -> mm_interconnect_0:Nios_V_data_manager_awprot
	wire  [31:0] nios_v_data_manager_wdata;                             // Nios_V:data_manager_wdata -> mm_interconnect_0:Nios_V_data_manager_wdata
	wire         nios_v_data_manager_arvalid;                           // Nios_V:data_manager_arvalid -> mm_interconnect_0:Nios_V_data_manager_arvalid
	wire         nios_v_data_manager_bvalid;                            // mm_interconnect_0:Nios_V_data_manager_bvalid -> Nios_V:data_manager_bvalid
	wire         nios_v_data_manager_awvalid;                           // Nios_V:data_manager_awvalid -> mm_interconnect_0:Nios_V_data_manager_awvalid
	wire         nios_v_data_manager_rvalid;                            // mm_interconnect_0:Nios_V_data_manager_rvalid -> Nios_V:data_manager_rvalid
	wire  [31:0] nios_v_instruction_manager_awaddr;                     // Nios_V:instruction_manager_awaddr -> mm_interconnect_0:Nios_V_instruction_manager_awaddr
	wire   [1:0] nios_v_instruction_manager_bresp;                      // mm_interconnect_0:Nios_V_instruction_manager_bresp -> Nios_V:instruction_manager_bresp
	wire         nios_v_instruction_manager_arready;                    // mm_interconnect_0:Nios_V_instruction_manager_arready -> Nios_V:instruction_manager_arready
	wire  [31:0] nios_v_instruction_manager_rdata;                      // mm_interconnect_0:Nios_V_instruction_manager_rdata -> Nios_V:instruction_manager_rdata
	wire   [3:0] nios_v_instruction_manager_wstrb;                      // Nios_V:instruction_manager_wstrb -> mm_interconnect_0:Nios_V_instruction_manager_wstrb
	wire         nios_v_instruction_manager_wready;                     // mm_interconnect_0:Nios_V_instruction_manager_wready -> Nios_V:instruction_manager_wready
	wire         nios_v_instruction_manager_awready;                    // mm_interconnect_0:Nios_V_instruction_manager_awready -> Nios_V:instruction_manager_awready
	wire         nios_v_instruction_manager_rready;                     // Nios_V:instruction_manager_rready -> mm_interconnect_0:Nios_V_instruction_manager_rready
	wire         nios_v_instruction_manager_bready;                     // Nios_V:instruction_manager_bready -> mm_interconnect_0:Nios_V_instruction_manager_bready
	wire         nios_v_instruction_manager_wvalid;                     // Nios_V:instruction_manager_wvalid -> mm_interconnect_0:Nios_V_instruction_manager_wvalid
	wire  [31:0] nios_v_instruction_manager_araddr;                     // Nios_V:instruction_manager_araddr -> mm_interconnect_0:Nios_V_instruction_manager_araddr
	wire   [2:0] nios_v_instruction_manager_arprot;                     // Nios_V:instruction_manager_arprot -> mm_interconnect_0:Nios_V_instruction_manager_arprot
	wire   [1:0] nios_v_instruction_manager_rresp;                      // mm_interconnect_0:Nios_V_instruction_manager_rresp -> Nios_V:instruction_manager_rresp
	wire   [2:0] nios_v_instruction_manager_awprot;                     // Nios_V:instruction_manager_awprot -> mm_interconnect_0:Nios_V_instruction_manager_awprot
	wire  [31:0] nios_v_instruction_manager_wdata;                      // Nios_V:instruction_manager_wdata -> mm_interconnect_0:Nios_V_instruction_manager_wdata
	wire         nios_v_instruction_manager_arvalid;                    // Nios_V:instruction_manager_arvalid -> mm_interconnect_0:Nios_V_instruction_manager_arvalid
	wire         nios_v_instruction_manager_bvalid;                     // mm_interconnect_0:Nios_V_instruction_manager_bvalid -> Nios_V:instruction_manager_bvalid
	wire         nios_v_instruction_manager_awvalid;                    // Nios_V:instruction_manager_awvalid -> mm_interconnect_0:Nios_V_instruction_manager_awvalid
	wire         nios_v_instruction_manager_rvalid;                     // mm_interconnect_0:Nios_V_instruction_manager_rvalid -> Nios_V:instruction_manager_rvalid
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;  // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;    // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest; // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;     // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;        // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;       // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;   // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_nios_v_dm_agent_readdata;            // Nios_V:dm_agent_readdata -> mm_interconnect_0:Nios_V_dm_agent_readdata
	wire         mm_interconnect_0_nios_v_dm_agent_waitrequest;         // Nios_V:dm_agent_waitrequest -> mm_interconnect_0:Nios_V_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_nios_v_dm_agent_address;             // mm_interconnect_0:Nios_V_dm_agent_address -> Nios_V:dm_agent_address
	wire         mm_interconnect_0_nios_v_dm_agent_read;                // mm_interconnect_0:Nios_V_dm_agent_read -> Nios_V:dm_agent_read
	wire         mm_interconnect_0_nios_v_dm_agent_readdatavalid;       // Nios_V:dm_agent_readdatavalid -> mm_interconnect_0:Nios_V_dm_agent_readdatavalid
	wire         mm_interconnect_0_nios_v_dm_agent_write;               // mm_interconnect_0:Nios_V_dm_agent_write -> Nios_V:dm_agent_write
	wire  [31:0] mm_interconnect_0_nios_v_dm_agent_writedata;           // mm_interconnect_0:Nios_V_dm_agent_writedata -> Nios_V:dm_agent_writedata
	wire  [31:0] mm_interconnect_0_nios_v_timer_sw_agent_readdata;      // Nios_V:timer_sw_agent_readdata -> mm_interconnect_0:Nios_V_timer_sw_agent_readdata
	wire         mm_interconnect_0_nios_v_timer_sw_agent_waitrequest;   // Nios_V:timer_sw_agent_waitrequest -> mm_interconnect_0:Nios_V_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_nios_v_timer_sw_agent_address;       // mm_interconnect_0:Nios_V_timer_sw_agent_address -> Nios_V:timer_sw_agent_address
	wire         mm_interconnect_0_nios_v_timer_sw_agent_read;          // mm_interconnect_0:Nios_V_timer_sw_agent_read -> Nios_V:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_nios_v_timer_sw_agent_byteenable;    // mm_interconnect_0:Nios_V_timer_sw_agent_byteenable -> Nios_V:timer_sw_agent_byteenable
	wire         mm_interconnect_0_nios_v_timer_sw_agent_readdatavalid; // Nios_V:timer_sw_agent_readdatavalid -> mm_interconnect_0:Nios_V_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_nios_v_timer_sw_agent_write;         // mm_interconnect_0:Nios_V_timer_sw_agent_write -> Nios_V:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_nios_v_timer_sw_agent_writedata;     // mm_interconnect_0:Nios_V_timer_sw_agent_writedata -> Nios_V:timer_sw_agent_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                  // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                    // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire  [14:0] mm_interconnect_0_sram_s1_address;                     // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                  // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                       // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                   // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                       // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         irq_mapper_receiver0_irq;                              // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire  [15:0] nios_v_platform_irq_rx_irq;                            // irq_mapper:sender_irq -> Nios_V:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [DEBUG:rst_n, mm_interconnect_0:DEBUG_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                    // rst_controller_001:reset_out -> [Nios_V:ndm_reset_in_reset, Nios_V:reset_reset, SRAM:reset, irq_mapper:reset, mm_interconnect_0:Nios_V_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                // rst_controller_001:reset_req -> [SRAM:reset_req, rst_translator:reset_req_in]

	altera_avalon_jtag_uart #(
		.readBufferDepth            (64),
		.readIRQThreshold           (8),
		.useRegistersForReadBuffer  (0),
		.useRegistersForWriteBuffer (0),
		.writeBufferDepth           (64),
		.writeIRQThreshold          (8),
		.printingMethod             (0),
		.FIFO_WIDTH                 (8),
		.WR_WIDTHU                  (6),
		.RD_WIDTHU                  (6),
		.write_le                   ("ON"),
		.read_le                    ("ON"),
		.HEX_WRITE_DEPTH_STR        (64),
		.HEX_READ_DEPTH_STR         (64),
		.legacySignalAllow          (0)
	) debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	Nios_V_Nios_V nios_v (
		.clk                          (clk_clk),                                               //                 clk.clk
		.reset_reset                  (rst_controller_001_reset_out_reset),                    //               reset.reset
		.platform_irq_rx_irq          (nios_v_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.ndm_reset_in_reset           (rst_controller_001_reset_out_reset),                    //        ndm_reset_in.reset
		.timer_sw_agent_address       (mm_interconnect_0_nios_v_timer_sw_agent_address),       //      timer_sw_agent.address
		.timer_sw_agent_byteenable    (mm_interconnect_0_nios_v_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_read          (mm_interconnect_0_nios_v_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_nios_v_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_write         (mm_interconnect_0_nios_v_timer_sw_agent_write),         //                    .write
		.timer_sw_agent_writedata     (mm_interconnect_0_nios_v_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_waitrequest   (mm_interconnect_0_nios_v_timer_sw_agent_waitrequest),   //                    .waitrequest
		.timer_sw_agent_readdatavalid (mm_interconnect_0_nios_v_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.instruction_manager_awaddr   (nios_v_instruction_manager_awaddr),                     // instruction_manager.awaddr
		.instruction_manager_awprot   (nios_v_instruction_manager_awprot),                     //                    .awprot
		.instruction_manager_awvalid  (nios_v_instruction_manager_awvalid),                    //                    .awvalid
		.instruction_manager_awready  (nios_v_instruction_manager_awready),                    //                    .awready
		.instruction_manager_wdata    (nios_v_instruction_manager_wdata),                      //                    .wdata
		.instruction_manager_wstrb    (nios_v_instruction_manager_wstrb),                      //                    .wstrb
		.instruction_manager_wvalid   (nios_v_instruction_manager_wvalid),                     //                    .wvalid
		.instruction_manager_wready   (nios_v_instruction_manager_wready),                     //                    .wready
		.instruction_manager_bresp    (nios_v_instruction_manager_bresp),                      //                    .bresp
		.instruction_manager_bvalid   (nios_v_instruction_manager_bvalid),                     //                    .bvalid
		.instruction_manager_bready   (nios_v_instruction_manager_bready),                     //                    .bready
		.instruction_manager_araddr   (nios_v_instruction_manager_araddr),                     //                    .araddr
		.instruction_manager_arprot   (nios_v_instruction_manager_arprot),                     //                    .arprot
		.instruction_manager_arvalid  (nios_v_instruction_manager_arvalid),                    //                    .arvalid
		.instruction_manager_arready  (nios_v_instruction_manager_arready),                    //                    .arready
		.instruction_manager_rdata    (nios_v_instruction_manager_rdata),                      //                    .rdata
		.instruction_manager_rresp    (nios_v_instruction_manager_rresp),                      //                    .rresp
		.instruction_manager_rvalid   (nios_v_instruction_manager_rvalid),                     //                    .rvalid
		.instruction_manager_rready   (nios_v_instruction_manager_rready),                     //                    .rready
		.data_manager_awaddr          (nios_v_data_manager_awaddr),                            //        data_manager.awaddr
		.data_manager_awprot          (nios_v_data_manager_awprot),                            //                    .awprot
		.data_manager_awvalid         (nios_v_data_manager_awvalid),                           //                    .awvalid
		.data_manager_awready         (nios_v_data_manager_awready),                           //                    .awready
		.data_manager_wdata           (nios_v_data_manager_wdata),                             //                    .wdata
		.data_manager_wstrb           (nios_v_data_manager_wstrb),                             //                    .wstrb
		.data_manager_wvalid          (nios_v_data_manager_wvalid),                            //                    .wvalid
		.data_manager_wready          (nios_v_data_manager_wready),                            //                    .wready
		.data_manager_bresp           (nios_v_data_manager_bresp),                             //                    .bresp
		.data_manager_bvalid          (nios_v_data_manager_bvalid),                            //                    .bvalid
		.data_manager_bready          (nios_v_data_manager_bready),                            //                    .bready
		.data_manager_araddr          (nios_v_data_manager_araddr),                            //                    .araddr
		.data_manager_arprot          (nios_v_data_manager_arprot),                            //                    .arprot
		.data_manager_arvalid         (nios_v_data_manager_arvalid),                           //                    .arvalid
		.data_manager_arready         (nios_v_data_manager_arready),                           //                    .arready
		.data_manager_rdata           (nios_v_data_manager_rdata),                             //                    .rdata
		.data_manager_rresp           (nios_v_data_manager_rresp),                             //                    .rresp
		.data_manager_rvalid          (nios_v_data_manager_rvalid),                            //                    .rvalid
		.data_manager_rready          (nios_v_data_manager_rready),                            //                    .rready
		.dm_agent_address             (mm_interconnect_0_nios_v_dm_agent_address),             //            dm_agent.address
		.dm_agent_read                (mm_interconnect_0_nios_v_dm_agent_read),                //                    .read
		.dm_agent_readdata            (mm_interconnect_0_nios_v_dm_agent_readdata),            //                    .readdata
		.dm_agent_write               (mm_interconnect_0_nios_v_dm_agent_write),               //                    .write
		.dm_agent_writedata           (mm_interconnect_0_nios_v_dm_agent_writedata),           //                    .writedata
		.dm_agent_waitrequest         (mm_interconnect_0_nios_v_dm_agent_waitrequest),         //                    .waitrequest
		.dm_agent_readdatavalid       (mm_interconnect_0_nios_v_dm_agent_readdatavalid),       //                    .readdatavalid
		.dbg_reset_out_reset          (nios_v_dbg_reset_out_reset)                             //       dbg_reset_out.reset
	);

	Nios_V_SRAM sram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),        //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	Nios_V_mm_interconnect_0 mm_interconnect_0 (
		.Nios_V_data_manager_awaddr               (nios_v_data_manager_awaddr),                            //                Nios_V_data_manager.awaddr
		.Nios_V_data_manager_awprot               (nios_v_data_manager_awprot),                            //                                   .awprot
		.Nios_V_data_manager_awvalid              (nios_v_data_manager_awvalid),                           //                                   .awvalid
		.Nios_V_data_manager_awready              (nios_v_data_manager_awready),                           //                                   .awready
		.Nios_V_data_manager_wdata                (nios_v_data_manager_wdata),                             //                                   .wdata
		.Nios_V_data_manager_wstrb                (nios_v_data_manager_wstrb),                             //                                   .wstrb
		.Nios_V_data_manager_wvalid               (nios_v_data_manager_wvalid),                            //                                   .wvalid
		.Nios_V_data_manager_wready               (nios_v_data_manager_wready),                            //                                   .wready
		.Nios_V_data_manager_bresp                (nios_v_data_manager_bresp),                             //                                   .bresp
		.Nios_V_data_manager_bvalid               (nios_v_data_manager_bvalid),                            //                                   .bvalid
		.Nios_V_data_manager_bready               (nios_v_data_manager_bready),                            //                                   .bready
		.Nios_V_data_manager_araddr               (nios_v_data_manager_araddr),                            //                                   .araddr
		.Nios_V_data_manager_arprot               (nios_v_data_manager_arprot),                            //                                   .arprot
		.Nios_V_data_manager_arvalid              (nios_v_data_manager_arvalid),                           //                                   .arvalid
		.Nios_V_data_manager_arready              (nios_v_data_manager_arready),                           //                                   .arready
		.Nios_V_data_manager_rdata                (nios_v_data_manager_rdata),                             //                                   .rdata
		.Nios_V_data_manager_rresp                (nios_v_data_manager_rresp),                             //                                   .rresp
		.Nios_V_data_manager_rvalid               (nios_v_data_manager_rvalid),                            //                                   .rvalid
		.Nios_V_data_manager_rready               (nios_v_data_manager_rready),                            //                                   .rready
		.Nios_V_instruction_manager_awaddr        (nios_v_instruction_manager_awaddr),                     //         Nios_V_instruction_manager.awaddr
		.Nios_V_instruction_manager_awprot        (nios_v_instruction_manager_awprot),                     //                                   .awprot
		.Nios_V_instruction_manager_awvalid       (nios_v_instruction_manager_awvalid),                    //                                   .awvalid
		.Nios_V_instruction_manager_awready       (nios_v_instruction_manager_awready),                    //                                   .awready
		.Nios_V_instruction_manager_wdata         (nios_v_instruction_manager_wdata),                      //                                   .wdata
		.Nios_V_instruction_manager_wstrb         (nios_v_instruction_manager_wstrb),                      //                                   .wstrb
		.Nios_V_instruction_manager_wvalid        (nios_v_instruction_manager_wvalid),                     //                                   .wvalid
		.Nios_V_instruction_manager_wready        (nios_v_instruction_manager_wready),                     //                                   .wready
		.Nios_V_instruction_manager_bresp         (nios_v_instruction_manager_bresp),                      //                                   .bresp
		.Nios_V_instruction_manager_bvalid        (nios_v_instruction_manager_bvalid),                     //                                   .bvalid
		.Nios_V_instruction_manager_bready        (nios_v_instruction_manager_bready),                     //                                   .bready
		.Nios_V_instruction_manager_araddr        (nios_v_instruction_manager_araddr),                     //                                   .araddr
		.Nios_V_instruction_manager_arprot        (nios_v_instruction_manager_arprot),                     //                                   .arprot
		.Nios_V_instruction_manager_arvalid       (nios_v_instruction_manager_arvalid),                    //                                   .arvalid
		.Nios_V_instruction_manager_arready       (nios_v_instruction_manager_arready),                    //                                   .arready
		.Nios_V_instruction_manager_rdata         (nios_v_instruction_manager_rdata),                      //                                   .rdata
		.Nios_V_instruction_manager_rresp         (nios_v_instruction_manager_rresp),                      //                                   .rresp
		.Nios_V_instruction_manager_rvalid        (nios_v_instruction_manager_rvalid),                     //                                   .rvalid
		.Nios_V_instruction_manager_rready        (nios_v_instruction_manager_rready),                     //                                   .rready
		.clk_0_clk_clk                            (clk_clk),                                               //                          clk_0_clk.clk
		.DEBUG_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                        //  DEBUG_reset_reset_bridge_in_reset.reset
		.Nios_V_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // Nios_V_reset_reset_bridge_in_reset.reset
		.DEBUG_avalon_jtag_slave_address          (mm_interconnect_0_debug_avalon_jtag_slave_address),     //            DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write            (mm_interconnect_0_debug_avalon_jtag_slave_write),       //                                   .write
		.DEBUG_avalon_jtag_slave_read             (mm_interconnect_0_debug_avalon_jtag_slave_read),        //                                   .read
		.DEBUG_avalon_jtag_slave_readdata         (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                                   .readdata
		.DEBUG_avalon_jtag_slave_writedata        (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                                   .writedata
		.DEBUG_avalon_jtag_slave_waitrequest      (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect       (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.Nios_V_dm_agent_address                  (mm_interconnect_0_nios_v_dm_agent_address),             //                    Nios_V_dm_agent.address
		.Nios_V_dm_agent_write                    (mm_interconnect_0_nios_v_dm_agent_write),               //                                   .write
		.Nios_V_dm_agent_read                     (mm_interconnect_0_nios_v_dm_agent_read),                //                                   .read
		.Nios_V_dm_agent_readdata                 (mm_interconnect_0_nios_v_dm_agent_readdata),            //                                   .readdata
		.Nios_V_dm_agent_writedata                (mm_interconnect_0_nios_v_dm_agent_writedata),           //                                   .writedata
		.Nios_V_dm_agent_readdatavalid            (mm_interconnect_0_nios_v_dm_agent_readdatavalid),       //                                   .readdatavalid
		.Nios_V_dm_agent_waitrequest              (mm_interconnect_0_nios_v_dm_agent_waitrequest),         //                                   .waitrequest
		.Nios_V_timer_sw_agent_address            (mm_interconnect_0_nios_v_timer_sw_agent_address),       //              Nios_V_timer_sw_agent.address
		.Nios_V_timer_sw_agent_write              (mm_interconnect_0_nios_v_timer_sw_agent_write),         //                                   .write
		.Nios_V_timer_sw_agent_read               (mm_interconnect_0_nios_v_timer_sw_agent_read),          //                                   .read
		.Nios_V_timer_sw_agent_readdata           (mm_interconnect_0_nios_v_timer_sw_agent_readdata),      //                                   .readdata
		.Nios_V_timer_sw_agent_writedata          (mm_interconnect_0_nios_v_timer_sw_agent_writedata),     //                                   .writedata
		.Nios_V_timer_sw_agent_byteenable         (mm_interconnect_0_nios_v_timer_sw_agent_byteenable),    //                                   .byteenable
		.Nios_V_timer_sw_agent_readdatavalid      (mm_interconnect_0_nios_v_timer_sw_agent_readdatavalid), //                                   .readdatavalid
		.Nios_V_timer_sw_agent_waitrequest        (mm_interconnect_0_nios_v_timer_sw_agent_waitrequest),   //                                   .waitrequest
		.SRAM_s1_address                          (mm_interconnect_0_sram_s1_address),                     //                            SRAM_s1.address
		.SRAM_s1_write                            (mm_interconnect_0_sram_s1_write),                       //                                   .write
		.SRAM_s1_readdata                         (mm_interconnect_0_sram_s1_readdata),                    //                                   .readdata
		.SRAM_s1_writedata                        (mm_interconnect_0_sram_s1_writedata),                   //                                   .writedata
		.SRAM_s1_byteenable                       (mm_interconnect_0_sram_s1_byteenable),                  //                                   .byteenable
		.SRAM_s1_chipselect                       (mm_interconnect_0_sram_s1_chipselect),                  //                                   .chipselect
		.SRAM_s1_clken                            (mm_interconnect_0_sram_s1_clken)                        //                                   .clken
	);

	Nios_V_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios_v_platform_irq_rx_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios_v_dbg_reset_out_reset),     // reset_in0.reset
		.reset_in1      (nios_v_dbg_reset_out_reset),     // reset_in1.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios_v_dbg_reset_out_reset),             // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
